module top_tb();

   initial begin
      $display("Hi");
   end

endmodule : top_tb
