module top_tb();

   TinyORAMCore oram(

		     );

   initial begin
      $display("Hi");
   end

endmodule : top_tb
